--STD_LOGIC >> for single bit 

a: STD_LOGIC; >> means>> the bit value could be 1,0,z(floating),...
a<= "1";

--STD_LOGIC_VICTOR >> for single bit 

a: STD_LOGIC_VICTOR(3 downto 0);>> means>>[3,2,1,0]  >> each single bit can contain 1,0,z(floating),...
a<= "1010";

0 >>means>> grounded 
1 >>means>> high
z >>means>> floating